`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Dimitris Christodoulou
// 
// Create Date:    15:04:14 11/21/2018 
// Design Name: 
// Module Name:    mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mem(RESET, CLK, ADDR, read_mem, read_mem_vertical, DO_RED, DO_GREEN, DO_BLUE);
input RESET, CLK, read_mem;
input read_mem_vertical;
input [13:0] ADDR;
output reg DO_RED, DO_GREEN, DO_BLUE;

wire red, green, blue;

	RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//RED 6 ROWS OF PIXEL
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//RED 6 ROWS OF PIXEL
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_0C(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_0D(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_0E(256'h00000000000000000000000000000000_00000000000000000000000000000000),//GREEN 6 ROWS OF PIXEL
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_12(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_13(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_14(256'h00000000000000000000000000000000_00000000000000000000000000000000),//GREEN 6 ROWS OF PIXEL
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_18(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_19(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1A(256'h00000000000000000000000000000000_00000000000000000000000000000000),//BLUE 6 ROWS OF PIXEL
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_1E(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1F(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000_00000000000000000000000000000000),//BLUE 6 ROWS OF PIXEL
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_24(256'h0F000F000F000F000F000F000F000F00_0F000F000F000F000F000F000F000F00),
      .INIT_25(256'h0F000F000F000F000F000F000F000F00_0F000F000F000F000F000F000F000F00),
      .INIT_26(256'h0F000F000F000F000F000F000F000F00_0F000F000F000F000F000F000F000F00),//BLACK SPACE (BLACK - RED - GREEN - BLUE)
      .INIT_27(256'hFF00FF00FF00FF00FF00FF00FF00FF00_FF00FF00FF00FF00FF00FF00FF00FF00),
      .INIT_28(256'hFF00FF00FF00FF00FF00FF00FF00FF00_FF00FF00FF00FF00FF00FF00FF00FF00),
      .INIT_29(256'hFF00FF00FF00FF00FF00FF00FF00FF00_FF00FF00FF00FF00FF00FF00FF00FF00),//WHITE SPACE (WHITE - RED - GREEN - BLUE)
      .INIT_2A(256'h0F000F000F000F000F000F000F000F00_0F000F000F000F000F000F000F000F00),
      .INIT_2B(256'h0F000F000F000F000F000F000F000F00_0F000F000F000F000F000F000F000F00),
      .INIT_2C(256'h0F000F000F000F000F000F000F000F00_0F000F000F000F000F000F000F000F00),//BLACK SPACE (BLACK - RED - GREEN - BLUE)
      .INIT_2D(256'hFF00FF00FF00FF00FF00FF00FF00FF00_FF00FF00FF00FF00FF00FF00FF00FF00),
      .INIT_2E(256'hFF00FF00FF00FF00FF00FF00FF00FF00_FF00FF00FF00FF00FF00FF00FF00FF00),
      .INIT_2F(256'hFF00FF00FF00FF00FF00FF00FF00FF00_FF00FF00FF00FF00FF00FF00FF00FF00),//WHITE SPACE (WHITE - RED - GREEN - BLUE)
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_red_inst (
      .DO(red),      // 1-bit Data Output
      .ADDR(ADDR),  // 14-bit Address Input
      .CLK(CLK),    // Clock
      .EN(1'b1),      // RAM Enable Input
      .SSR(RESET),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );
	
	
	RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_01(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_02(256'h00000000000000000000000000000000_00000000000000000000000000000000),//RED 6 ROWS OF PIXEL
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_06(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_07(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_08(256'h00000000000000000000000000000000_00000000000000000000000000000000),//RED 6 ROWS OF PIXEL
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//GREEN 6 ROWS OF PIXEL
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//GREEN 6 ROWS OF PIXEL
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_18(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_19(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1A(256'h00000000000000000000000000000000_00000000000000000000000000000000),//BLUE 6 ROWS OF PIXEL
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_1E(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1F(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000_00000000000000000000000000000000),//BLUE 6 ROWS OF PIXEL
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_24(256'h00F000F000F000F000F000F000F000F0_00F000F000F000F000F000F000F000F0),
      .INIT_25(256'h00F000F000F000F000F000F000F000F0_00F000F000F000F000F000F000F000F0),
      .INIT_26(256'h00F000F000F000F000F000F000F000F0_00F000F000F000F000F000F000F000F0),//BLACK SPACE (BLACK - RED - GREEN - BLUE)
      .INIT_27(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0_F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),
      .INIT_28(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0_F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),
      .INIT_29(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0_F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),//WHITE SPACE (WHITE - RED - GREEN - BLUE)
      .INIT_2A(256'h00F000F000F000F000F000F000F000F0_00F000F000F000F000F000F000F000F0),
      .INIT_2B(256'h00F000F000F000F000F000F000F000F0_00F000F000F000F000F000F000F000F0),
      .INIT_2C(256'h00F000F000F000F000F000F000F000F0_00F000F000F000F000F000F000F000F0),//BLACK SPACE (BLACK - RED - GREEN - BLUE)
      .INIT_2D(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0_F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),
      .INIT_2E(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0_F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),
      .INIT_2F(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0_F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),//WHITE SPACE (WHITE - RED - GREEN - BLUE)
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_green_inst (
      .DO(green),      // 1-bit Data Output
      .ADDR(ADDR),  // 14-bit Address Input
      .CLK(CLK),    // Clock
      .EN(1'b1),      // RAM Enable Input
      .SSR(RESET),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );
	
	
	RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_01(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_02(256'h00000000000000000000000000000000_00000000000000000000000000000000),//RED 6 ROWS OF PIXEL
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_06(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_07(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_08(256'h00000000000000000000000000000000_00000000000000000000000000000000),//RED 6 ROWS OF PIXEL
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_0C(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_0D(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_0E(256'h00000000000000000000000000000000_00000000000000000000000000000000),//GREEN 6 ROWS OF PIXEL
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_12(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_13(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_14(256'h00000000000000000000000000000000_00000000000000000000000000000000),//GREEN 6 ROWS OF PIXEL
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//BLUE 6 ROWS OF PIXEL
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 8192 to 12287
      .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//BLUE 6 ROWS OF PIXEL
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//WHITE 6 ROWS OF PIXEL
      .INIT_24(256'h000F000F000F000F000F000F000F000F_000F000F000F000F000F000F000F000F),
      .INIT_25(256'h000F000F000F000F000F000F000F000F_000F000F000F000F000F000F000F000F),
      .INIT_26(256'h000F000F000F000F000F000F000F000F_000F000F000F000F000F000F000F000F),//BLACK SPACE (RED - GREEN - BLUE - BLACK - BLACK)
      .INIT_27(256'hF00FF00FF00FF00FF00FF00FF00FF00F_F00FF00FF00FF00FF00FF00FF00FF00F),
      .INIT_28(256'hF00FF00FF00FF00FF00FF00FF00FF00F_F00FF00FF00FF00FF00FF00FF00FF00F),
      .INIT_29(256'hF00FF00FF00FF00FF00FF00FF00FF00F_F00FF00FF00FF00FF00FF00FF00FF00F),//WHITE SPACE (WHITE - RED - GREEN - BLUE)
      .INIT_2A(256'h000F000F000F000F000F000F000F000F_000F000F000F000F000F000F000F000F),
      .INIT_2B(256'h000F000F000F000F000F000F000F000F_000F000F000F000F000F000F000F000F),
      .INIT_2C(256'h000F000F000F000F000F000F000F000F_000F000F000F000F000F000F000F000F),//BLACK SPACE (RED - GREEN - BLUE - BLACK - BLACK)
      .INIT_2D(256'hF00FF00FF00FF00FF00FF00FF00FF00F_F00FF00FF00FF00FF00FF00FF00FF00F),
      .INIT_2E(256'hF00FF00FF00FF00FF00FF00FF00FF00F_F00FF00FF00FF00FF00FF00FF00FF00F),
      .INIT_2F(256'hF00FF00FF00FF00FF00FF00FF00FF00F_F00FF00FF00FF00FF00FF00FF00FF00F),//WHITE SPACE (WHITE - RED - GREEN - BLUE)
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_blue_inst (
      .DO(blue),      // 1-bit Data Output
      .ADDR(ADDR),  // 14-bit Address Input
      .CLK(CLK),    // Clock
      .EN(1'b1),      // RAM Enable Input
      .SSR(RESET),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );
	
	always@(posedge CLK or posedge RESET)
	begin
		if(RESET)
		begin
			DO_RED = 1'b0;
			DO_GREEN = 1'b0;
			DO_BLUE = 1'b0;
		end
		else
		begin
			if(read_mem && read_mem_vertical)
			begin
				DO_RED = red;
				DO_GREEN = green;
				DO_BLUE = blue;
			end
			else
			begin
				DO_RED = 1'b0;
				DO_GREEN = 1'b0;
				DO_BLUE = 1'b0;
			end
		end
	end

endmodule
